interface out_b_if(input logic clk);

    logic out_valid_b;
    logic out_ready_b;
    logic [31:0]  out_instr_b;

endinterface
