interface out_a_if(input logic clk);

    logic out_valid_a;
    logic out_ready_a;
    logic [31:0]  out_instr_a;

endinterface
