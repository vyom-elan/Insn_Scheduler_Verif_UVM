interface out_d_if(input logic clk);

    logic out_valid_d;
    logic out_ready_d;
    logic [31:0]  out_instr_d;

endinterface
