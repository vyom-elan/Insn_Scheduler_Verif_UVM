interface out_c_if(input logic clk);

    logic out_valid_c;
    logic out_ready_c;
    logic [31:0]  out_instr_c;

endinterface
